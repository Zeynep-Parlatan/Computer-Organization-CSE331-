module my_and(
	input [31:0] first,
	input [31:0] second,
	output [31:0] result
);


and a0(result[31], first[31], second[31]);
and a1(result[30], first[30], second[30]);
and a2(result[29], first[29], second[29]);
and a3(result[28], first[28], second[28]);
and a4(result[27], first[27], second[27]);
and a5(result[26], first[26], second[26]);
and a6(result[25], first[25], second[25]);
and a7(result[24], first[24], second[24]);
and a8(result[23], first[23], second[23]);
and a9(result[22], first[22], second[22]);
and a10(result[21], first[21], second[21]);
and a11(result[20], first[20], second[20]);
and a12(result[19], first[19], second[19]);
and a13(result[18], first[18], second[18]);
and a14(result[17], first[17], second[17]);
and a15(result[16], first[16], second[16]);
and a16(result[15], first[15], second[15]);
and a17(result[14], first[14], second[14]);
and a18(result[13], first[13], second[13]);
and a19(result[12], first[12], second[12]);
and a20(result[11], first[11], second[11]);
and a21(result[10], first[10], second[10]);
and a22(result[9], first[9], second[9]);
and a23(result[8], first[8], second[8]);
and a24(result[7], first[7], second[7]);
and a25(result[6], first[6], second[6]);
and a26(result[5], first[5], second[5]);
and a27(result[4], first[4], second[4]);
and a28(result[3], first[3], second[3]);
and a29(result[2], first[2], second[2]);
and a30(result[1], first[1], second[1]);
and a31(result[0], first[0], second[0]);

endmodule
